library verilog;
use verilog.vl_types.all;
entity diplay_tester_vlg_vec_tst is
end diplay_tester_vlg_vec_tst;
